library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

package data_package is
  
  type DATA_ARRAY is array ( 2 downto 0) of signed( 15 downto 0);
  
end data_package;