--**************************************************************************************************
--
--  
--
--**************************************************************************************************
--  Comprehensive VHDL                  
--  Mumma Radar Lab                 
--  Hamdi Abdelbagi                 
--  ALU TB
--   9/18/2016
--**************************************************************************************************
--
--  
--
--**************************************************************************************************



entity ALU_TB is
end;

library IEEE;
use IEEE.Std_logic_1164.all;
use IEEE.Numeric_Std.all;

architecture Bench of ALU_TB is

  constant OP_SIZE       : POSITIVE := 4;

  -- Signals connected to the ALU
  signal Cout, Equal : Std_logic;
  signal F: std_logic_vector(7 downto 0);
  signal A, B: std_logic_vector(7 downto 0) := (others => '0');
  signal Op: std_logic_vector(OP_SIZE-1 downto 0);

  -- Some interesting values for A and B. The test
  -- assigns every combination of these to A and B
  -- for each operation
  constant Value0: Std_logic_vector := "00000000";
  constant Value1: Std_logic_vector := "00000001";
  constant Value2: Std_logic_vector := "00000011";
  constant Value3: Std_logic_vector := "00001000";
  constant Value4: Std_logic_vector := "00001111";
  constant Value5: Std_logic_vector := "10000000";
  constant Value6: Std_logic_vector := "11111000";
  constant Value7: Std_logic_vector := "11111111";

  constant NUM_VALUES    : POSITIVE := 8;
  constant NUM_OP_VALUES : POSITIVE := 2 ** OP_SIZE;
  constant NUM_VECTORS   : POSITIVE := NUM_VALUES * NUM_VALUES * NUM_OP_VALUES;

  -- Delay constants
  constant OP_DELAY : TIME := 10 ns;
  constant  A_DELAY : TIME := NUM_OP_VALUES * OP_DELAY;
  constant  B_DELAY : TIME := NUM_VALUES * A_DELAY;

  -- Expected result and error recording
  signal Exp : Std_logic_vector(1 to 10);
  constant DONT_CARE : Std_logic_vector(7 downto 0) := "--------";

  signal     F_Error_count : NATURAL := 0;
  signal  Cout_Error_count : NATURAL := 0;
  signal Equal_Error_count : NATURAL := 0;

  signal     F_OK : BOOLEAN := TRUE;
  signal  Cout_OK : BOOLEAN := TRUE;
  signal Equal_OK : BOOLEAN := TRUE;

begin

  UUT: entity WORK.ALU(A1)
    port map ( A     => A,
               B     => B,
               Op    => Op,
               F     => F,
               Cout  => Cout,
               Equal => Equal);

  -- Assigns B once to each test value
  BStim: process
  begin
    B <= Value0;
    wait for B_DELAY;
    B <= Value1;
    wait for B_DELAY;
    B <= Value2;
    wait for B_DELAY;
    B <= Value3;
    wait for B_DELAY;
    B <= Value4;
    wait for B_DELAY;
    B <= Value5;
    wait for B_DELAY;
    B <= Value6;
    wait for B_DELAY;
    B <= Value7;
    wait for B_DELAY;
    wait;
  end process BStim;

  -- Assigns A to each test value in turn
  -- for each different value of B
  AStim: process
  begin
    for I in 1 to NUM_VALUES loop
      A <= Value0;
      wait for A_DELAY;
      A <= Value1;
      wait for A_DELAY;
      A <= Value2;
      wait for A_DELAY;
      A <= Value3;
      wait for A_DELAY;
      A <= Value4;
      wait for A_DELAY;
      A <= Value5;
      wait for A_DELAY;
      A <= Value6;
      wait for A_DELAY;
      A <= Value7;
      wait for A_DELAY;
    end loop;
    wait;
  end process AStim;

  -- Assigns Op to each possible value (including the
  -- unused ones) for every combination of A and B
  OpStim: process
  begin
    for I in 1 to NUM_VALUES * NUM_VALUES loop
      for J in 0 to NUM_OP_VALUES-1 loop
        Op <= Std_logic_vector(To_unsigned(J,4));
        wait for OP_DELAY;
      end loop;
    end loop;
    wait;
  end process OpStim;

  -- Assigned the expected output values to "Exp".
  Expected: process
  begin
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000001001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000101"; wait for OP_DELAY;
    Exp <= "0000000101"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0000001001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000001001"; wait for OP_DELAY;
    Exp <= "1000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100100"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000111000"; wait for OP_DELAY;
    Exp <= "1111001010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000110"; wait for OP_DELAY;
    Exp <= "0111111110"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "1111011110"; wait for OP_DELAY;
    Exp <= "0000100100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000011001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000001101"; wait for OP_DELAY;
    Exp <= "0000001101"; wait for OP_DELAY;
    Exp <= "1111110111"; wait for OP_DELAY;
    Exp <= "1111110111"; wait for OP_DELAY;
    Exp <= "0000011001"; wait for OP_DELAY;
    Exp <= "0000000101"; wait for OP_DELAY;
    Exp <= "0000011001"; wait for OP_DELAY;
    Exp <= "1000000101"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0000101100"; wait for OP_DELAY;
    Exp <= "0000010100"; wait for OP_DELAY;
    Exp <= "1111101110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001001000"; wait for OP_DELAY;
    Exp <= "0000110000"; wait for OP_DELAY;
    Exp <= "1111010010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000001110"; wait for OP_DELAY;
    Exp <= "0111110110"; wait for OP_DELAY;
    Exp <= "1000001100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111101110"; wait for OP_DELAY;
    Exp <= "1111010110"; wait for OP_DELAY;
    Exp <= "0000101100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1111110010"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100100"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000101100"; wait for OP_DELAY;
    Exp <= "1111101110"; wait for OP_DELAY;
    Exp <= "0000010100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000100001"; wait for OP_DELAY;
    Exp <= "0000100001"; wait for OP_DELAY;
    Exp <= "1111100011"; wait for OP_DELAY;
    Exp <= "1111100011"; wait for OP_DELAY;
    Exp <= "0001000001"; wait for OP_DELAY;
    Exp <= "0000010001"; wait for OP_DELAY;
    Exp <= "0001000001"; wait for OP_DELAY;
    Exp <= "0000010001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0001011100"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000100010"; wait for OP_DELAY;
    Exp <= "0111100010"; wait for OP_DELAY;
    Exp <= "1000100000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "1111011110"; wait for OP_DELAY;
    Exp <= "0000100100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "1111001010"; wait for OP_DELAY;
    Exp <= "0000111000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001001000"; wait for OP_DELAY;
    Exp <= "1111010010"; wait for OP_DELAY;
    Exp <= "0000110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001011100"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0001111001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000111101"; wait for OP_DELAY;
    Exp <= "0000111101"; wait for OP_DELAY;
    Exp <= "1111000111"; wait for OP_DELAY;
    Exp <= "1111000111"; wait for OP_DELAY;
    Exp <= "0001111001"; wait for OP_DELAY;
    Exp <= "0000011101"; wait for OP_DELAY;
    Exp <= "0001111001"; wait for OP_DELAY;
    Exp <= "1000011101"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "1000111110"; wait for OP_DELAY;
    Exp <= "0111000110"; wait for OP_DELAY;
    Exp <= "1000111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "1110100110"; wait for OP_DELAY;
    Exp <= "0001011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000111000"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000110"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "0111111110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000001110"; wait for OP_DELAY;
    Exp <= "1000001100"; wait for OP_DELAY;
    Exp <= "0111110110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000100010"; wait for OP_DELAY;
    Exp <= "1000100000"; wait for OP_DELAY;
    Exp <= "0111100010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000111110"; wait for OP_DELAY;
    Exp <= "1000111100"; wait for OP_DELAY;
    Exp <= "0111000110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000011"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "1000000011"; wait for OP_DELAY;
    Exp <= "1000000011"; wait for OP_DELAY;
    Exp <= "1000000001"; wait for OP_DELAY;
    Exp <= "1000000001"; wait for OP_DELAY;
    Exp <= "0000000011"; wait for OP_DELAY;
    Exp <= "0100000001"; wait for OP_DELAY;
    Exp <= "0000000111"; wait for OP_DELAY;
    Exp <= "0100000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0111100010"; wait for OP_DELAY;
    Exp <= "0111100000"; wait for OP_DELAY;
    Exp <= "1000100010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0111111110"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1000000110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "0000100100"; wait for OP_DELAY;
    Exp <= "1111011110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111101110"; wait for OP_DELAY;
    Exp <= "0000101100"; wait for OP_DELAY;
    Exp <= "1111010110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001011100"; wait for OP_DELAY;
    Exp <= "1110100110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0111100010"; wait for OP_DELAY;
    Exp <= "1000100010"; wait for OP_DELAY;
    Exp <= "0111100000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111000011"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "1111100011"; wait for OP_DELAY;
    Exp <= "1111100011"; wait for OP_DELAY;
    Exp <= "0000100001"; wait for OP_DELAY;
    Exp <= "0000100001"; wait for OP_DELAY;
    Exp <= "1111000011"; wait for OP_DELAY;
    Exp <= "0111110001"; wait for OP_DELAY;
    Exp <= "1111000111"; wait for OP_DELAY;
    Exp <= "0111110001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "1111011110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1111111010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000001000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "1111110010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000001100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111110110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000011000"; wait for OP_DELAY;
    Exp <= "1000000100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0000100100"; wait for OP_DELAY;
    Exp <= "1111011110"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "0000010000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000111000"; wait for OP_DELAY;
    Exp <= "0001000000"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000111100"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "0001111000"; wait for OP_DELAY;
    Exp <= "1000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0111111110"; wait for OP_DELAY;
    Exp <= "1000000110"; wait for OP_DELAY;
    Exp <= "0111111100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1000000010"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1000000000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "0000000010"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "0000000110"; wait for OP_DELAY;
    Exp <= "0100000000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111011110"; wait for OP_DELAY;
    Exp <= "1111100110"; wait for OP_DELAY;
    Exp <= "0000011100"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "1111100010"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "0000100000"; wait for OP_DELAY;
    Exp <= "0000000100"; wait for OP_DELAY;
    Exp <= "1111000010"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "1111000110"; wait for OP_DELAY;
    Exp <= "0111110000"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "---------0"; wait for OP_DELAY;
    Exp <= "0000000000"; wait for OP_DELAY;
    Exp <= "1111111110"; wait for OP_DELAY;
    Exp <= "1111111011"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "0000000101"; wait for OP_DELAY;
    Exp <= "0000000101"; wait for OP_DELAY;
    Exp <= "1111111011"; wait for OP_DELAY;
    Exp <= "0111111101"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    Exp <= "1111111101"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "---------1"; wait for OP_DELAY;
    Exp <= "0000000001"; wait for OP_DELAY;
    Exp <= "1111111111"; wait for OP_DELAY;
    wait;
  end process Expected;

  -- Checks the outputs are as expected. An expected "don't care"
  -- value ('-') means the corresponding output is ignored.
  Check : process
  begin
    wait for OP_DELAY - 1 NS;
    for I in 1 to NUM_VECTORS loop
      if ( Exp(1 to 8) /= DONT_CARE ) and ( F /= Exp(1 to 8) ) then
        F_OK              <= FALSE;
        F_Error_count     <= F_Error_Count + 1;
      end if;
      if ( Exp(9) /= '-' ) and ( Cout /= Exp(9) ) then
        Cout_OK           <= FALSE;
        Cout_Error_count  <= Cout_Error_Count + 1;
      end if;
      if ( Exp(10) /= '-' ) and ( Equal /= Exp(10) ) then
        Equal_OK          <= FALSE;
        Equal_Error_count <= Equal_Error_Count + 1;
      end if;
      wait for OP_DELAY;
    end loop;
    
    if F_Error_count = 0 and Cout_Error_count = 0 and 
       Equal_error_count = 0 then
       report "ALU Finished OK";
    else
       report "ALU Finished with ERRORS";
    end if;
    wait;
  end process Check;

end architecture Bench;
